----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:24:06 01/13/2025 
-- Design Name: 
-- Module Name:    RAM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity RAM is
    Port (
        i_clk : in std_logic;
        i_en_a : in std_logic;
        i_addr_a : in std_logic_vector (11 downto 0);
        i_we_a : in std_logic_vector (3 downto 0);
        i_data_a : in std_logic_vector (31 downto 0);
        o_data_a : out std_logic_vector (31 downto 0);
        i_clk_b : in std_logic;
        i_en_b : in std_logic;
        i_addr_b : in std_logic_vector (11 downto 0);
        i_we_b : in std_logic_vector (3 downto 0);
        i_data_b : in std_logic_vector (31 downto 0);
        o_data_b : out std_logic_vector (31 downto 0)
    );
end RAM;

architecture Behavioral of RAM is

    signal s_addr_a : std_logic_vector(13 downto 0) := (others => '0');
    signal s_addr_b : std_logic_vector(13 downto 0) := (others => '0');
    
    signal s_en_a : std_logic_vector(7 downto 0) := (others => '0');
    signal s_en_b : std_logic_vector(7 downto 0) := (others => '0');
    
    signal s_o_data_a_0 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_a_1 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_a_2 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_a_3 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_a_4 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_a_5 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_a_6 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_a_7 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_b_0 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_b_1 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_b_2 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_b_3 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_b_4 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_b_5 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_b_6 : std_logic_vector(31 downto 0) := (others => '0');
    signal s_o_data_b_7 : std_logic_vector(31 downto 0) := (others => '0');

begin

    RAMB16BWER_inst_0 : RAMB16BWER
    generic map (
        -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
        DATA_WIDTH_A => 36,
        DATA_WIDTH_B => 36,
        -- DOA_REG/DOB_REG: Optional output register (0 or 1)
        DOA_REG => 0,
        DOB_REG => 0,
        -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
        EN_RSTRAM_A => TRUE,
        EN_RSTRAM_B => TRUE,
        -- INITP_00 to INITP_07: Initial memory contents.
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INIT_00 to INIT_3F: Initial memory contents.
        INIT_00 => X"018555130007A503200007B70000006F161000EF2C8000EF0001011300010117",
        INIT_01 => X"02C798630100031300C886930088871300000793200008B70000806700157513",
        INIT_02 => X"2006661300A7202303F67613FFF60613FE079CE30027F7930007278320000737",
        INIT_03 => X"0105883300279813FE081CE3008878130008A8030000806700C7A223200007B7",
        INIT_04 => X"0027F7930007278320000737FADFF06F0066A023010720230017879300082803",
        INIT_05 => X"0006851300E6A22324076713200006B703F77713FFF6071300A72023FE079CE3",
        INIT_06 => X"0027969300072803FE069CE30206F693000526830000806700C7946300868713",
        INIT_07 => X"11312E231321202312912223ED010113FD9FF06F001787930106A02300D586B3",
        INIT_08 => X"FE050EE3EFDFF0EF00060913000584930005099311412C231281242312112623",
        INIT_09 => X"20000A3700C12623000405930009851306961463000006130004079301010413",
        INIT_0A => X"000405930009851300C12603020792631007F793FFE00513000A2783EE9FF0EF",
        INIT_0B => X"124124831281240312C12083040782632007F793FFD00513000A2783F35FF0EF",
        INIT_0C => X"00478793001606130127A023000080671301011311812A0311C1298312012903",
        INIT_0D => X"FB9FF06F00000513FE9798E30017879301271A630044041300042703F8DFF06F",
        INIT_0E => X"BF0585930331262300001437000015B702812C23FC010113FB1FF06FFFF00513",
        INIT_0F => X"02112E2301812C2301712E23036120230351222302912A23C884051300050993",
        INIT_10 => X"01000C1302000A9300001BB700001B3771C000EF000004930341242303212823",
        INIT_11 => X"C884051300C10593158000EF0FF4F51300C10593700000EFC8840513C2CB0593",
        INIT_12 => X"012A07B30000091301498A336D8000EF00449A13C8840513C30B85936E8000EF",
        INIT_13 => X"020005936B0000EFC884051300C10593120000EF0019091300C105930007C503",
        INIT_14 => X"F95492E3660000EF00148493C884051300A00593FD891AE3674000EFC8840513",
        INIT_15 => X"02012B0302412A8302812A0302C1298303012903034124830381240303C12083",
        INIT_16 => X"009122230000143700812423FF010113000080670401011301812C0301C12B83",
        INIT_17 => X"004124830081240300C1208300F46C63C9048793000014B7C8C4041300112623",
        INIT_18 => X"02812423FD010113FD9FF06F000780E700440413000427830000806701010113",
        INIT_19 => X"0211262300C10513C4458593000504930110061302912223000015B700058413",
        INIT_1A => X"002787B30207879300F7F79340E4D7B3FFC0061301C0071300040693788000EF",
        INIT_1B => X"0281240302C1208300040423FEC710E3FEF68FA300168693FFC70713FEC7C783",
        INIT_1C => X"02812423000015B70005849302912223FD010113000080670301011302412483",
        INIT_1D => X"0207879300445793714000EF0211262300C10513C44585930005041301100613",
        INIT_1E => X"FEC44783002784330204079300F480230004812300F47413FEC7C783002787B3",
        INIT_1F => X"00B52023000502230000806703010113024124830281240302C1208300F480A3",
        INIT_20 => X"004547830000806700B7802300B502230005278300F5E5B30045478300008067",
        INIT_21 => X"00C5222300B520230000806700B7802300B502230005278300F5F5B30015B593",
        INIT_22 => X"FA9FF06F0010059300452503FCDFF06F00100593004525030000806700D52423",
        INIT_23 => X"0004A503FDDFF0EF00A0041300050493001126230091222300812423FF010113",
        INIT_24 => X"004124830081240300C12083FE0416E3330000EF0FF474130FF00593FFF40413",
        INIT_25 => X"000604930005041300912A2300812C2300112E23FE0101130000806701010113",
        INIT_26 => X"2E0000EF0FF0059300042503F85FF0EF00058993000689130131262301212823",
        INIT_27 => X"2C0000EF0184D593000425032CC000EF0409E59300042503F65FF0EF00040513",
        INIT_28 => X"2A0000EF0FF5F5930084D593000425032B0000EF0FF5F5930104D59300042503",
        INIT_29 => X"280000EF0FF009130019659300042503290000EF008004930FF4F59300042503",
        INIT_2A => X"0181240301C12083FE0496E3FFF4849301251663274000EF0FF0059300042503",
        INIT_2B => X"0005049300912223FF010113000080670201011300C129830101290301412483",
        INIT_2C => X"0004A50300050413228000EF0121202300812423001126230FF0059300052503",
        INIT_2D => X"200000EF0FF005930004A50300A4643301051513214000EF018414130FF00593",
        INIT_2E => X"008124030085653300C120831EC000EF008919130FF005930004A50300050913",
        INIT_2F => X"0081242300112623FF01011300008067010101130001290300A9653300412483",
        INIT_30 => X"E8DFF0EF00040513000005930000061309400693E59FF0EF0005041300912223",
        INIT_31 => X"08A7E6630005049300100793E79FF0EF00040513008005931AA0061308600693",
        INIT_32 => X"00040513E51FF0EF0004051303A005930000061300000693F31FF0EF00040513",
        INIT_33 => X"4000063700000693E35FF0EF00040513037005930000061300000693F15FF0EF",
        INIT_34 => X"28C000EFC5858593000015B700842503FC051CE3E21FF0EF0004051302900593",
        INIT_35 => X"EB9FF0EF0004051300050493DF9FF0EF0004051303A005930000061300000693",
        INIT_36 => X"000080670101011300412483000485130081240300C12083D91FF0EF00040513",
        INIT_37 => X"0006049300058913000504130121282300912A2300812C2300112E23FE010113",
        INIT_38 => X"0FF00793D91FF0EF00040513011005930000069300090613D45FF0EF01312623",
        INIT_39 => X"080000EF0FF005930004250300078993387909130000193706F5046300050913",
        INIT_3A => X"0FF005930004250320048913FE0912E30109591301091913FFF9091301351A63",
        INIT_3B => X"040000EF0FE009130FF0059300042503FE9916E3FEA48FA3058000EF00148493",
        INIT_3C => X"014124830181240301C12083CC5FF0EF00040513034000EF0FF0059300042503",
        INIT_3D => X"000527030000806700B520230000806702010113010129030009051300C12983",
        INIT_3E => X"FE078CE30047F793001747830005270300B70023FE078CE30047F79300174783",
        INIT_3F => X"00B780A30005278300008067003575130017C503000527830000806700074503",
        -- INIT_A/INIT_B: Initial values on output port
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- INIT_FILE: Optional file used to specify initial RAM contents
        INIT_FILE => "NONE",
        -- RSTTYPE: "SYNC" or "ASYNC" 
        RSTTYPE => "SYNC",
        -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
        RST_PRIORITY_A => "CE",
        RST_PRIORITY_B => "CE",
        -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
        SIM_COLLISION_CHECK => "ALL",
        -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
        SIM_DEVICE => "SPARTAN6",
        -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        WRITE_MODE_A => "WRITE_FIRST",
        WRITE_MODE_B => "WRITE_FIRST" 
    )
    port map (
        -- Port A Data: 32-bit (each) output: Port A data
        DOA => s_o_data_a_0,       -- 32-bit output: A port data output
        DOPA => open,     -- 4-bit output: A port parity output
        -- Port B Data: 32-bit (each) output: Port B data
        DOB => s_o_data_b_0,       -- 32-bit output: B port data output
        DOPB => open,     -- 4-bit output: B port parity output
        -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
        ADDRA => s_addr_a,   -- 14-bit input: A port address input
        CLKA => i_clk,     -- 1-bit input: A port clock input
        ENA => s_en_a(0),       -- 1-bit input: A port enable input
        REGCEA => '1', -- 1-bit input: A port register clock enable input
        RSTA => '0',     -- 1-bit input: A port register set/reset input
        WEA => i_we_a,       -- 4-bit input: Port A byte-wide write enable input
        -- Port A Data: 32-bit (each) input: Port A data
        DIA => i_data_a,       -- 32-bit input: A port data input
        DIPA => "0000",     -- 4-bit input: A port parity input
        -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
        ADDRB => s_addr_b,   -- 14-bit input: B port address input
        CLKB => i_clk_b,     -- 1-bit input: B port clock input
        ENB => s_en_b(0),       -- 1-bit input: B port enable input
        REGCEB => '1', -- 1-bit input: B port register clock enable input
        RSTB => '0',     -- 1-bit input: B port register set/reset input
        WEB => i_we_b,       -- 4-bit input: Port B byte-wide write enable input
        -- Port B Data: 32-bit (each) input: Port B data
        DIB => i_data_b,       -- 32-bit input: B port data input
        DIPB => "0000"      -- 4-bit input: B port parity input
    );
    
    RAMB16BWER_inst_1 : RAMB16BWER
    generic map (
        -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
        DATA_WIDTH_A => 36,
        DATA_WIDTH_B => 36,
        -- DOA_REG/DOB_REG: Optional output register (0 or 1)
        DOA_REG => 0,
        DOB_REG => 0,
        -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
        EN_RSTRAM_A => TRUE,
        EN_RSTRAM_B => TRUE,
        -- INITP_00 to INITP_07: Initial memory contents.
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INIT_00 to INIT_3F: Initial memory contents.
        INIT_00 => X"001005130000806700A035330027C503000718630037C7030005278300008067",
        INIT_01 => X"0000806700B781230005278300E781A30FF5F5930085D7130005278300008067",
        INIT_02 => X"0006A5030007A58300052683004527830000806700B522230045859300B52023",
        INIT_03 => X"00149413008124230005849300912223FF01011300008067FEE59AE30007A703",
        INIT_04 => X"FB5FF0EF00050913001126230024141301212023009404330034141300940433",
        INIT_05 => X"FE9568E300B41463FE85ECE3FA1FF0EF0009051300B404330084B43300A404B3",
        INIT_06 => X"40B787B300559793000080670101011300012903004124830081240300C12083",
        INIT_07 => X"00174783000527030000806700B52023F81FF06F0035959300B785B300279793",
        INIT_08 => X"FE079CE30027F79300174783000527030000806700B70023FE079CE30047F793",
        INIT_09 => X"0005841300050493001126230091222300812423FF0101130000806700074503",
        INIT_0A => X"000485130000806701010113004124830081240300C1208300059C6300044583",
        INIT_0B => X"20112623C845051307C00593DF01011300001537FD9FF06F00140413F99FF0EF",
        INIT_0C => X"000015B7F41FF0EFC6C405133E800593E99FF0EF000014372091222320812423",
        INIT_0D => X"00010613C3DFF0EFC6048513000014B7F7DFF0EFC8850513C385859300001537",
        INIT_0E => X"000106131C6155831C815783FF8FF0EF00010513D19FF0EFC604851300000593",
        INIT_0F => X"C7448513000014B7FD4FF0EF00010513CF5FF0EFC604851300B7E5B301079793",
        INIT_10 => X"A01FF0EF00100593C7448513EC9FF0EF1F400593C6C40513A01FF0EF00100593",
        INIT_11 => X"C88905130000193701212023FF010113FD1FF06FEB1FF0EFC6C405131F400593",
        INIT_12 => X"C8440513100005B700001437EA1FF0EF009122230081242300112623100005B7",
        INIT_13 => X"00001537981FF0EF00458593C7C48513100025B7000014B7D51FF0EF01058593",
        INIT_14 => X"C6050513C7C48613C8890693C844059300001537971FF0EFC7450513100025B7",
        INIT_15 => X"C6C50513100015B700001537000129030041248300C1208300812403999FF0EF",
        INIT_16 => X"06C7F263003007930607966300C508B30037F79300A5C7B3D7DFF06F01010113",
        INIT_17 => X"0005869306D7C4630200079340E606B3FFC8F6130C079A630005071300357793",
        INIT_18 => X"FFF60613FEC7E8E3FF07AE2300468693004787930006A80302C77A6300070793",
        INIT_19 => X"000080670117686300C7073300C585B30047071300458593FFC6761340E60633",
        INIT_1A => X"00008067FEE898E3FEF70FA300158593001707130005C783FF157CE300050713",
        INIT_1B => X"0185A3030145AE030105AE8300C5AF030085AF830045A2830005A3830205A683",
        INIT_1C => X"FFE72423FFF72223FE57202340E606B3FC772E23FED72E230247071301C5A803",
        INIT_1D => X"0005C683F45FF06FFAD7C6E302458593FF072C23FE672A23FFC72823FFD72623",
        INIT_1E => X"00377793001707130005C683F0078EE300158593FED70FA30037779300170713",
        INIT_1F => X"32302031302030302020202020202020F01FF06FFC079AE300158593FED70FA3",
        INIT_20 => X"3020433020423020413020393020383020373020363020353020343020333020",
        INIT_21 => X"7075207265776F500000000020203A2000007830000000000A46302045302044",
        INIT_22 => X"00000A796461655200000000464544434241393837363534333231300000000A",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000A30000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INIT_A/INIT_B: Initial values on output port
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- INIT_FILE: Optional file used to specify initial RAM contents
        INIT_FILE => "NONE",
        -- RSTTYPE: "SYNC" or "ASYNC" 
        RSTTYPE => "SYNC",
        -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
        RST_PRIORITY_A => "CE",
        RST_PRIORITY_B => "CE",
        -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
        SIM_COLLISION_CHECK => "ALL",
        -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
        SIM_DEVICE => "SPARTAN6",
        -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        WRITE_MODE_A => "WRITE_FIRST",
        WRITE_MODE_B => "WRITE_FIRST" 
    )
    port map (
        -- Port A Data: 32-bit (each) output: Port A data
        DOA => s_o_data_a_1,       -- 32-bit output: A port data output
        DOPA => open,     -- 4-bit output: A port parity output
        -- Port B Data: 32-bit (each) output: Port B data
        DOB => s_o_data_b_1,       -- 32-bit output: B port data output
        DOPB => open,     -- 4-bit output: B port parity output
        -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
        ADDRA => s_addr_a,   -- 14-bit input: A port address input
        CLKA => i_clk,     -- 1-bit input: A port clock input
        ENA => s_en_a(1),       -- 1-bit input: A port enable input
        REGCEA => '1', -- 1-bit input: A port register clock enable input
        RSTA => '0',     -- 1-bit input: A port register set/reset input
        WEA => i_we_a,       -- 4-bit input: Port A byte-wide write enable input
        -- Port A Data: 32-bit (each) input: Port A data
        DIA => i_data_a,       -- 32-bit input: A port data input
        DIPA => "0000",     -- 4-bit input: A port parity input
        -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
        ADDRB => s_addr_b,   -- 14-bit input: B port address input
        CLKB => i_clk_b,     -- 1-bit input: B port clock input
        ENB => s_en_b(1),       -- 1-bit input: B port enable input
        REGCEB => '1', -- 1-bit input: B port register clock enable input
        RSTB => '0',     -- 1-bit input: B port register set/reset input
        WEB => i_we_b,       -- 4-bit input: Port B byte-wide write enable input
        -- Port B Data: 32-bit (each) input: Port B data
        DIB => i_data_b,       -- 32-bit input: B port data input
        DIPB => "0000"      -- 4-bit input: B port parity input
    );
    
    RAMB16BWER_inst_2 : RAMB16BWER
    generic map (
        -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
        DATA_WIDTH_A => 36,
        DATA_WIDTH_B => 36,
        -- DOA_REG/DOB_REG: Optional output register (0 or 1)
        DOA_REG => 0,
        DOB_REG => 0,
        -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
        EN_RSTRAM_A => TRUE,
        EN_RSTRAM_B => TRUE,
        -- INITP_00 to INITP_07: Initial memory contents.
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INIT_00 to INIT_3F: Initial memory contents.
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000022",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000", --32B
        -- INIT_A/INIT_B: Initial values on output port
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- INIT_FILE: Optional file used to specify initial RAM contents
        INIT_FILE => "NONE",
        -- RSTTYPE: "SYNC" or "ASYNC" 
        RSTTYPE => "SYNC",
        -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
        RST_PRIORITY_A => "CE",
        RST_PRIORITY_B => "CE",
        -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
        SIM_COLLISION_CHECK => "ALL",
        -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
        SIM_DEVICE => "SPARTAN6",
        -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        WRITE_MODE_A => "WRITE_FIRST",
        WRITE_MODE_B => "WRITE_FIRST" 
    )
    port map (
        -- Port A Data: 32-bit (each) output: Port A data
        DOA => s_o_data_a_2,       -- 32-bit output: A port data output
        DOPA => open,     -- 4-bit output: A port parity output
        -- Port B Data: 32-bit (each) output: Port B data
        DOB => s_o_data_b_2,       -- 32-bit output: B port data output
        DOPB => open,     -- 4-bit output: B port parity output
        -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
        ADDRA => s_addr_a,   -- 14-bit input: A port address input
        CLKA => i_clk,     -- 1-bit input: A port clock input
        ENA => s_en_a(2),       -- 1-bit input: A port enable input
        REGCEA => '1', -- 1-bit input: A port register clock enable input
        RSTA => '0',     -- 1-bit input: A port register set/reset input
        WEA => i_we_a,       -- 4-bit input: Port A byte-wide write enable input
        -- Port A Data: 32-bit (each) input: Port A data
        DIA => i_data_a,       -- 32-bit input: A port data input
        DIPA => "0000",     -- 4-bit input: A port parity input
        -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
        ADDRB => s_addr_b,   -- 14-bit input: B port address input
        CLKB => i_clk_b,     -- 1-bit input: B port clock input
        ENB => s_en_b(2),       -- 1-bit input: B port enable input
        REGCEB => '1', -- 1-bit input: B port register clock enable input
        RSTB => '0',     -- 1-bit input: B port register set/reset input
        WEB => i_we_b,       -- 4-bit input: Port B byte-wide write enable input
        -- Port B Data: 32-bit (each) input: Port B data
        DIB => i_data_b,       -- 32-bit input: B port data input
        DIPB => "0000"      -- 4-bit input: B port parity input
    );
    
    RAMB16BWER_inst_3 : RAMB16BWER
    generic map (
        -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
        DATA_WIDTH_A => 36,
        DATA_WIDTH_B => 36,
        -- DOA_REG/DOB_REG: Optional output register (0 or 1)
        DOA_REG => 0,
        DOB_REG => 0,
        -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
        EN_RSTRAM_A => TRUE,
        EN_RSTRAM_B => TRUE,
        -- INITP_00 to INITP_07: Initial memory contents.
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INIT_00 to INIT_3F: Initial memory contents.
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000033",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000", --32B
        -- INIT_A/INIT_B: Initial values on output port
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- INIT_FILE: Optional file used to specify initial RAM contents
        INIT_FILE => "NONE",
        -- RSTTYPE: "SYNC" or "ASYNC" 
        RSTTYPE => "SYNC",
        -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
        RST_PRIORITY_A => "CE",
        RST_PRIORITY_B => "CE",
        -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
        SIM_COLLISION_CHECK => "ALL",
        -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
        SIM_DEVICE => "SPARTAN6",
        -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        WRITE_MODE_A => "WRITE_FIRST",
        WRITE_MODE_B => "WRITE_FIRST" 
    )
    port map (
        -- Port A Data: 32-bit (each) output: Port A data
        DOA => s_o_data_a_3,       -- 32-bit output: A port data output
        DOPA => open,     -- 4-bit output: A port parity output
        -- Port B Data: 32-bit (each) output: Port B data
        DOB => s_o_data_b_3,       -- 32-bit output: B port data output
        DOPB => open,     -- 4-bit output: B port parity output
        -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
        ADDRA => s_addr_a,   -- 14-bit input: A port address input
        CLKA => i_clk,     -- 1-bit input: A port clock input
        ENA => s_en_a(3),       -- 1-bit input: A port enable input
        REGCEA => '1', -- 1-bit input: A port register clock enable input
        RSTA => '0',     -- 1-bit input: A port register set/reset input
        WEA => i_we_a,       -- 4-bit input: Port A byte-wide write enable input
        -- Port A Data: 32-bit (each) input: Port A data
        DIA => i_data_a,       -- 32-bit input: A port data input
        DIPA => "0000",     -- 4-bit input: A port parity input
        -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
        ADDRB => s_addr_b,   -- 14-bit input: B port address input
        CLKB => i_clk_b,     -- 1-bit input: B port clock input
        ENB => s_en_b(3),       -- 1-bit input: B port enable input
        REGCEB => '1', -- 1-bit input: B port register clock enable input
        RSTB => '0',     -- 1-bit input: B port register set/reset input
        WEB => i_we_b,       -- 4-bit input: Port B byte-wide write enable input
        -- Port B Data: 32-bit (each) input: Port B data
        DIB => i_data_b,       -- 32-bit input: B port data input
        DIPB => "0000"      -- 4-bit input: B port parity input
    );
    
    RAMB16BWER_inst_4 : RAMB16BWER
    generic map (
        -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
        DATA_WIDTH_A => 36,
        DATA_WIDTH_B => 36,
        -- DOA_REG/DOB_REG: Optional output register (0 or 1)
        DOA_REG => 0,
        DOB_REG => 0,
        -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
        EN_RSTRAM_A => TRUE,
        EN_RSTRAM_B => TRUE,
        -- INITP_00 to INITP_07: Initial memory contents.
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INIT_00 to INIT_3F: Initial memory contents.
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000044",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000", --32B
        -- INIT_A/INIT_B: Initial values on output port
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- INIT_FILE: Optional file used to specify initial RAM contents
        INIT_FILE => "NONE",
        -- RSTTYPE: "SYNC" or "ASYNC" 
        RSTTYPE => "SYNC",
        -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
        RST_PRIORITY_A => "CE",
        RST_PRIORITY_B => "CE",
        -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
        SIM_COLLISION_CHECK => "ALL",
        -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
        SIM_DEVICE => "SPARTAN6",
        -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        WRITE_MODE_A => "WRITE_FIRST",
        WRITE_MODE_B => "WRITE_FIRST" 
    )
    port map (
        -- Port A Data: 32-bit (each) output: Port A data
        DOA => s_o_data_a_4,       -- 32-bit output: A port data output
        DOPA => open,     -- 4-bit output: A port parity output
        -- Port B Data: 32-bit (each) output: Port B data
        DOB => s_o_data_b_4,       -- 32-bit output: B port data output
        DOPB => open,     -- 4-bit output: B port parity output
        -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
        ADDRA => s_addr_a,   -- 14-bit input: A port address input
        CLKA => i_clk,     -- 1-bit input: A port clock input
        ENA => s_en_a(4),       -- 1-bit input: A port enable input
        REGCEA => '1', -- 1-bit input: A port register clock enable input
        RSTA => '0',     -- 1-bit input: A port register set/reset input
        WEA => i_we_a,       -- 4-bit input: Port A byte-wide write enable input
        -- Port A Data: 32-bit (each) input: Port A data
        DIA => i_data_a,       -- 32-bit input: A port data input
        DIPA => "0000",     -- 4-bit input: A port parity input
        -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
        ADDRB => s_addr_b,   -- 14-bit input: B port address input
        CLKB => i_clk_b,     -- 1-bit input: B port clock input
        ENB => s_en_b(4),       -- 1-bit input: B port enable input
        REGCEB => '1', -- 1-bit input: B port register clock enable input
        RSTB => '0',     -- 1-bit input: B port register set/reset input
        WEB => i_we_b,       -- 4-bit input: Port B byte-wide write enable input
        -- Port B Data: 32-bit (each) input: Port B data
        DIB => i_data_b,       -- 32-bit input: B port data input
        DIPB => "0000"      -- 4-bit input: B port parity input
    );
    
    RAMB16BWER_inst_5 : RAMB16BWER
    generic map (
        -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
        DATA_WIDTH_A => 36,
        DATA_WIDTH_B => 36,
        -- DOA_REG/DOB_REG: Optional output register (0 or 1)
        DOA_REG => 0,
        DOB_REG => 0,
        -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
        EN_RSTRAM_A => TRUE,
        EN_RSTRAM_B => TRUE,
        -- INITP_00 to INITP_07: Initial memory contents.
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INIT_00 to INIT_3F: Initial memory contents.
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000055",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000", --32B
        -- INIT_A/INIT_B: Initial values on output port
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- INIT_FILE: Optional file used to specify initial RAM contents
        INIT_FILE => "NONE",
        -- RSTTYPE: "SYNC" or "ASYNC" 
        RSTTYPE => "SYNC",
        -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
        RST_PRIORITY_A => "CE",
        RST_PRIORITY_B => "CE",
        -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
        SIM_COLLISION_CHECK => "ALL",
        -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
        SIM_DEVICE => "SPARTAN6",
        -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        WRITE_MODE_A => "WRITE_FIRST",
        WRITE_MODE_B => "WRITE_FIRST" 
    )
    port map (
        -- Port A Data: 32-bit (each) output: Port A data
        DOA => s_o_data_a_5,       -- 32-bit output: A port data output
        DOPA => open,     -- 4-bit output: A port parity output
        -- Port B Data: 32-bit (each) output: Port B data
        DOB => s_o_data_b_5,       -- 32-bit output: B port data output
        DOPB => open,     -- 4-bit output: B port parity output
        -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
        ADDRA => s_addr_a,   -- 14-bit input: A port address input
        CLKA => i_clk,     -- 1-bit input: A port clock input
        ENA => s_en_a(5),       -- 1-bit input: A port enable input
        REGCEA => '1', -- 1-bit input: A port register clock enable input
        RSTA => '0',     -- 1-bit input: A port register set/reset input
        WEA => i_we_a,       -- 4-bit input: Port A byte-wide write enable input
        -- Port A Data: 32-bit (each) input: Port A data
        DIA => i_data_a,       -- 32-bit input: A port data input
        DIPA => "0000",     -- 4-bit input: A port parity input
        -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
        ADDRB => s_addr_b,   -- 14-bit input: B port address input
        CLKB => i_clk_b,     -- 1-bit input: B port clock input
        ENB => s_en_b(5),       -- 1-bit input: B port enable input
        REGCEB => '1', -- 1-bit input: B port register clock enable input
        RSTB => '0',     -- 1-bit input: B port register set/reset input
        WEB => i_we_b,       -- 4-bit input: Port B byte-wide write enable input
        -- Port B Data: 32-bit (each) input: Port B data
        DIB => i_data_b,       -- 32-bit input: B port data input
        DIPB => "0000"      -- 4-bit input: B port parity input
    );
    
    RAMB16BWER_inst_6 : RAMB16BWER
    generic map (
        -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
        DATA_WIDTH_A => 36,
        DATA_WIDTH_B => 36,
        -- DOA_REG/DOB_REG: Optional output register (0 or 1)
        DOA_REG => 0,
        DOB_REG => 0,
        -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
        EN_RSTRAM_A => TRUE,
        EN_RSTRAM_B => TRUE,
        -- INITP_00 to INITP_07: Initial memory contents.
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INIT_00 to INIT_3F: Initial memory contents.
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000066",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000", --32B
        -- INIT_A/INIT_B: Initial values on output port
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- INIT_FILE: Optional file used to specify initial RAM contents
        INIT_FILE => "NONE",
        -- RSTTYPE: "SYNC" or "ASYNC" 
        RSTTYPE => "SYNC",
        -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
        RST_PRIORITY_A => "CE",
        RST_PRIORITY_B => "CE",
        -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
        SIM_COLLISION_CHECK => "ALL",
        -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
        SIM_DEVICE => "SPARTAN6",
        -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        WRITE_MODE_A => "WRITE_FIRST",
        WRITE_MODE_B => "WRITE_FIRST" 
    )
    port map (
        -- Port A Data: 32-bit (each) output: Port A data
        DOA => s_o_data_a_6,       -- 32-bit output: A port data output
        DOPA => open,     -- 4-bit output: A port parity output
        -- Port B Data: 32-bit (each) output: Port B data
        DOB => s_o_data_b_6,       -- 32-bit output: B port data output
        DOPB => open,     -- 4-bit output: B port parity output
        -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
        ADDRA => s_addr_a,   -- 14-bit input: A port address input
        CLKA => i_clk,     -- 1-bit input: A port clock input
        ENA => s_en_a(6),       -- 1-bit input: A port enable input
        REGCEA => '1', -- 1-bit input: A port register clock enable input
        RSTA => '0',     -- 1-bit input: A port register set/reset input
        WEA => i_we_a,       -- 4-bit input: Port A byte-wide write enable input
        -- Port A Data: 32-bit (each) input: Port A data
        DIA => i_data_a,       -- 32-bit input: A port data input
        DIPA => "0000",     -- 4-bit input: A port parity input
        -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
        ADDRB => s_addr_b,   -- 14-bit input: B port address input
        CLKB => i_clk_b,     -- 1-bit input: B port clock input
        ENB => s_en_b(6),       -- 1-bit input: B port enable input
        REGCEB => '1', -- 1-bit input: B port register clock enable input
        RSTB => '0',     -- 1-bit input: B port register set/reset input
        WEB => i_we_b,       -- 4-bit input: Port B byte-wide write enable input
        -- Port B Data: 32-bit (each) input: Port B data
        DIB => i_data_b,       -- 32-bit input: B port data input
        DIPB => "0000"      -- 4-bit input: B port parity input
    );
    
    RAMB16BWER_inst_7 : RAMB16BWER
    generic map (
        -- DATA_WIDTH_A/DATA_WIDTH_B: 0, 1, 2, 4, 9, 18, or 36
        DATA_WIDTH_A => 36,
        DATA_WIDTH_B => 36,
        -- DOA_REG/DOB_REG: Optional output register (0 or 1)
        DOA_REG => 0,
        DOB_REG => 0,
        -- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
        EN_RSTRAM_A => TRUE,
        EN_RSTRAM_B => TRUE,
        -- INITP_00 to INITP_07: Initial memory contents.
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INIT_00 to INIT_3F: Initial memory contents.
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000077",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000", --32B
        -- INIT_A/INIT_B: Initial values on output port
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- INIT_FILE: Optional file used to specify initial RAM contents
        INIT_FILE => "NONE",
        -- RSTTYPE: "SYNC" or "ASYNC" 
        RSTTYPE => "SYNC",
        -- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR" 
        RST_PRIORITY_A => "CE",
        RST_PRIORITY_B => "CE",
        -- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE" 
        SIM_COLLISION_CHECK => "ALL",
        -- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
        SIM_DEVICE => "SPARTAN6",
        -- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- WRITE_MODE_A/WRITE_MODE_B: "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        WRITE_MODE_A => "WRITE_FIRST",
        WRITE_MODE_B => "WRITE_FIRST" 
    )
    port map (
        -- Port A Data: 32-bit (each) output: Port A data
        DOA => s_o_data_a_7,       -- 32-bit output: A port data output
        DOPA => open,     -- 4-bit output: A port parity output
        -- Port B Data: 32-bit (each) output: Port B data
        DOB => s_o_data_b_7,       -- 32-bit output: B port data output
        DOPB => open,     -- 4-bit output: B port parity output
        -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals
        ADDRA => s_addr_a,   -- 14-bit input: A port address input
        CLKA => i_clk,     -- 1-bit input: A port clock input
        ENA => s_en_a(7),       -- 1-bit input: A port enable input
        REGCEA => '1', -- 1-bit input: A port register clock enable input
        RSTA => '0',     -- 1-bit input: A port register set/reset input
        WEA => i_we_a,       -- 4-bit input: Port A byte-wide write enable input
        -- Port A Data: 32-bit (each) input: Port A data
        DIA => i_data_a,       -- 32-bit input: A port data input
        DIPA => "0000",     -- 4-bit input: A port parity input
        -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals
        ADDRB => s_addr_b,   -- 14-bit input: B port address input
        CLKB => i_clk_b,     -- 1-bit input: B port clock input
        ENB => s_en_b(7),       -- 1-bit input: B port enable input
        REGCEB => '1', -- 1-bit input: B port register clock enable input
        RSTB => '0',     -- 1-bit input: B port register set/reset input
        WEB => i_we_b,       -- 4-bit input: Port B byte-wide write enable input
        -- Port B Data: 32-bit (each) input: Port B data
        DIB => i_data_b,       -- 32-bit input: B port data input
        DIPB => "0000"      -- 4-bit input: B port parity input
    );
    
    process(i_addr_a, i_en_a)
    begin
        case i_addr_a(11 downto 9) is
            when "000" =>
                s_en_a <= "0000000" & i_en_a;
            when "001" =>
                s_en_a <= "000000" & i_en_a & "0";
            when "010" =>
                s_en_a <= "00000" & i_en_a & "00";
            when "011" =>
                s_en_a <= "0000" & i_en_a & "000";
            when "100" =>
                s_en_a <= "000" & i_en_a & "0000";
            when "101" =>
                s_en_a <= "00" & i_en_a & "00000";
            when "110" =>
                s_en_a <= "0" & i_en_a & "000000";
            when "111" =>
                s_en_a <= i_en_a & "0000000";
            when others =>
                s_en_a <= (others => '0');
        end case;
    end process;
    
    process(i_addr_b, i_en_b)
    begin
        case i_addr_b(11 downto 9) is
            when "000" =>
                s_en_b <= "0000000" & i_en_b;
            when "001" =>
                s_en_b <= "000000" & i_en_b & "0";
            when "010" =>
                s_en_b <= "00000" & i_en_b & "00";
            when "011" =>
                s_en_b <= "0000" & i_en_b & "000";
            when "100" =>
                s_en_b <= "000" & i_en_b & "0000";
            when "101" =>
                s_en_b <= "00" & i_en_b & "00000";
            when "110" =>
                s_en_b <= "0" & i_en_b & "000000";
            when "111" =>
                s_en_b <= i_en_b & "0000000";
            when others =>
                s_en_b <= (others => '0');
        end case;
    end process;
    
    process(i_addr_a, s_o_data_a_0, s_o_data_a_1, s_o_data_a_2, s_o_data_a_3, s_o_data_a_4, s_o_data_a_5, s_o_data_a_6, s_o_data_a_7)
    begin
        case i_addr_a(11 downto 9) is
            when "000" =>
                o_data_a <= s_o_data_a_0;
            when "001" =>
                o_data_a <= s_o_data_a_1;
            when "010" =>
                o_data_a <= s_o_data_a_2;
            when "011" =>
                o_data_a <= s_o_data_a_3;
            when "100" =>
                o_data_a <= s_o_data_a_4;
            when "101" =>
                o_data_a <= s_o_data_a_5;
            when "110" =>
                o_data_a <= s_o_data_a_6;
            when "111" =>
                o_data_a <= s_o_data_a_7;
            when others =>
                o_data_a <= (others => '0');
        end case;
    end process;
    
    process(i_addr_b, s_o_data_b_0, s_o_data_b_1, s_o_data_b_2, s_o_data_b_3, s_o_data_b_4, s_o_data_b_5, s_o_data_b_6, s_o_data_b_7)
    begin
        case i_addr_b(11 downto 9) is
            when "000" =>
                o_data_b <= s_o_data_b_0;
            when "001" =>
                o_data_b <= s_o_data_b_1;
            when "010" =>
                o_data_b <= s_o_data_b_2;
            when "011" =>
                o_data_b <= s_o_data_b_3;
            when "100" =>
                o_data_b <= s_o_data_b_4;
            when "101" =>
                o_data_b <= s_o_data_b_5;
            when "110" =>
                o_data_b <= s_o_data_b_6;
            when "111" =>
                o_data_b <= s_o_data_b_7;
            when others =>
                o_data_b <= (others => '0');
        end case;
    end process;

    s_addr_a <= i_addr_a(8 downto 0) & "00000";
    s_addr_b <= i_addr_b(8 downto 0) & "00000";

end Behavioral;

